module ictest(A,B);
    input A;
    output B;
    assign B=A;
endmodule